//
// lab5a : version 08/13/2022
// 
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module sr_latch (output logic qa, output logic qb, input logic s,
	input logic r);

   // Enter your code here ...
   //
   assign qa = ~(s | qb);
   assign qb = ~(r | qa);

endmodule
