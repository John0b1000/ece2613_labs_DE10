// [Copy and paste the testbench template here]
