//
// lab5a : version 08/13/2022
// 
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module lvl_sen_sr_latch (output logic q, input logic s, input logic r,
	input logic c);
	
	// Enter your code here ...

endmodule
