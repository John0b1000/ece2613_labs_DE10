//
// lab6 : version 08/13/2022
// 
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module lab6_alu_1 (
	output logic c_out,
	output logic [6:0] cathode,
	input logic [11:0] sw
	);

	// Enter your code here ...

endmodule
