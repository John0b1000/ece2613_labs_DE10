//
// lab5a : version 08/13/2022
// 
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module d_flip_flop (output logic q, input logic d, input logic clk);

	// Enter your code here ...

endmodule
