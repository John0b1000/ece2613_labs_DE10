//
// lab7 : version 08/17/2022
//
`timescale 1ns / 1ps

module rotation_counter (output logic [6:0] cathode, output logic [3:0] anode,
	output logic error, input logic q_a, q_b, input logic rst, input logic clk);
	
	// Enter your code here ...

endmodule
