//
// lab2 : version 08/13/2022
// 
`timescale 1ns / 1ps
module hamming7_4_encode(
	output logic [7:1] e,
	input logic [4:1] d
	);

	// Enter your code here ...

endmodule
