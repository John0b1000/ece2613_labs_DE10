//
// lab3 : version 08/13/2022
//
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module lab3_decoder(
	output logic [3:0] an,
	output logic [6:0] cathode,
	input logic [6:0] sw
	);

	// Enter your code here ...

endmodule
