//
// lab5a : version 08/13/2022
// 
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
//////////////////////////////////////////////////////////////////////////////////
module transparent_d_latch (output logic q, input logic d, input logic c);

	// Enter your design here ...
	//
	lvl_sen_sr_latch u_lvl (.q(q), .s(d), .c(c), .r(~d));

endmodule
